module func_3 (
                input a,b,
                output func
              );
  and myAnd(func, a, b);
              
endmodule
