module func_2(
              input a,b,
              output func
            );

  assign func = a & b;            


endmodule
